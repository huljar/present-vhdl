library ieee;
use ieee.std_logic_1164.all;

entity sub_layer is
    port(data_in:  in std_logic_vector(63 downto 0);
         data_out: out std_logic_vector(63 downto 0)
    );
end sub_layer;

architecture behavioral of sub_layer is
    component sbox
        port(sbox_in:  in std_logic_vector(3 downto 0);
             sbox_out: out std_logic_vector(3 downto 0)
        );
    end component;

    begin
        GEN_SBOXES: for i in 15 downto 0 generate
            SX: sbox port map(
                sbox_in => data_in(4*i+3 downto 4*i),
                sbox_out => data_out(4*i+3 downto 4*i)
            );
        end generate;
    end behavioral;
